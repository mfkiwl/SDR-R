-- THIS IS A DUMMY FILE
-- NEED TO GENERATE A FIFO W/ XILINX IP
-- FIRST WORD FALL THRU ENABLED
-- 16 BITS INTO FIFO
--  8 BITS FROM FIFO
-- WILL DOCUMENT FURTHER
